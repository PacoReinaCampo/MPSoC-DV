`ifndef PERIPHERAL_UVM_DEFINES
`define PERIPHERAL_UVM_DEFINES

`define ADDER_WIDTH 4 
`define NO_OF_TRANSACTIONS 2000

`endif
