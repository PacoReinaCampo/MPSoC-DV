/*
 * Copyright 2018 Google LLC
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

package or1k_instr_test_pkg;

  import uvm_pkg::*;
  import or1k_instr_pkg::*;

  `include "or1k_instr_base_test.sv"
  `include "or1k_instr_test_lib.sv"
  `include "or1k_instr_cov_test.sv"

endpackage
