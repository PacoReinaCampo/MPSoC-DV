`define PERIPHERAL_UVM_KIT_VERSION "1.0ea"
`define PERIPHERAL_UVM_KIT_DATE "2010-04-30"
