`DEFINE_FC_INSTR(C_FLW,   CL_FORMAT, LOAD, OMSP32FC, UIMM)
`DEFINE_FC_INSTR(C_FSW,   CS_FORMAT, STORE, OMSP32FC, UIMM)
`DEFINE_FC_INSTR(C_FLWSP, CI_FORMAT, LOAD, OMSP32FC, UIMM)
`DEFINE_FC_INSTR(C_FSWSP, CSS_FORMAT, STORE, OMSP32FC, UIMM)
